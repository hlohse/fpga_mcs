
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity mcs_top is
  generic (
		hasDram: integer := 1;
		hasMbrot: integer := 0;
		xga: integer := 1; -- xga or 720p on hdmi
		hasHdmiTx: integer := 1;
		hasHdmiRx: integer := 0;
		simulation: integer := 0;
		trace: integer := 1;  -- use chipscope
    num_cx: integer := 800;
    num_mbpipe_stages: integer := 16
  );
  port (
		Clk : IN STD_LOGIC;
		Rst_n : IN STD_LOGIC;
		------------------------------------
		----- DRAM ports -------------------
		mcb3_dram_ck          : out std_logic;
		mcb3_dram_ck_n        : out std_logic;
		mcb3_dram_a           : out std_logic_vector(12 downto 0);
		mcb3_dram_ba          : out std_logic_vector(2 downto 0);
		mcb3_dram_ras_n       : out std_logic;
		mcb3_dram_cas_n       : out std_logic;
		mcb3_dram_we_n        : out std_logic;
		mcb3_dram_odt         : out std_logic;
		mcb3_dram_cke         : out std_logic;
		mcb3_dram_dq          : inout std_logic_vector(15 downto 0);
		mcb3_dram_dqs         : inout std_logic;
		mcb3_dram_dqs_n : inout std_logic;
		mcb3_dram_udqs   : inout std_logic;
		mcb3_dram_udm    : out std_logic; 
		mcb3_dram_udqs_n : inout std_logic;
		mcb3_dram_dm : out std_logic;
		mcb3_rzq                             : inout std_logic;
		mcb3_zio                              : inout std_logic;
		------------------------------------
		------ DRAM CS is not generated by MIG ---
		-- insert, if required (not on Atlys)
		-- mcb3_dram_cs_n        : out std_logic;
		--
		----- HDMI out ports ---------------
		hdmiTx0_p : OUT std_logic;
		hdmiTx0_n : OUT std_logic;
		hdmiTx1_p : OUT std_logic;
		hdmiTx1_n : OUT std_logic;
		hdmiTx2_p : OUT std_logic;
		hdmiTx2_n : OUT std_logic;
		hdmiTx3_p : OUT std_logic;
		hdmiTx3_n : OUT std_logic;
		------------------------------------
		------------------------------------
		UART_Rx : IN STD_LOGIC;
		UART_Tx : OUT STD_LOGIC;
		GPO1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		GPI1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		GPI2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    shiftPipe_debug: OUT STD_LOGIC_VECTOR(4 downto 0)
  );

end entity;
  
architecture rtl of mcs_top is

-- the core with trace option enabled
COMPONENT mblaze
  PORT (
    Clk : IN STD_LOGIC;
    Reset : IN STD_LOGIC;
    IO_Addr_Strobe : OUT STD_LOGIC;
    IO_Read_Strobe : OUT STD_LOGIC;
    IO_Write_Strobe : OUT STD_LOGIC;
    IO_Address : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    IO_Byte_Enable : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    IO_Write_Data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    IO_Read_Data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    IO_Ready : IN STD_LOGIC;
    UART_Rx : IN STD_LOGIC;
    UART_Tx : OUT STD_LOGIC;
    UART_Interrupt : OUT STD_LOGIC;
    FIT1_Interrupt : OUT STD_LOGIC;
    FIT1_Toggle : OUT STD_LOGIC;
    FIT2_Interrupt : OUT STD_LOGIC;
    FIT2_Toggle : OUT STD_LOGIC;
    PIT1_Interrupt : OUT STD_LOGIC;
    PIT1_Toggle : OUT STD_LOGIC;
    PIT2_Enable : IN STD_LOGIC;
    PIT2_Interrupt : OUT STD_LOGIC;
    PIT2_Toggle : OUT STD_LOGIC;
    GPO1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    GPI1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    GPI2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    GPI1_Interrupt : OUT STD_LOGIC;  -- GPI Interrupts are not enabled in MCS design
    GPI2_Interrupt : OUT STD_LOGIC;  -- GPI Interrupts are not enabled in MCS design
    INTC_Interrupt : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    INTC_IRQ : OUT STD_LOGIC;
    Trace_Instruction : OUT STD_LOGIC_VECTOR(0 TO 31);
    Trace_Valid_Instr : OUT STD_LOGIC;
    Trace_PC : OUT STD_LOGIC_VECTOR(0 TO 31);
    Trace_Reg_Write : OUT STD_LOGIC;
    Trace_Reg_Addr : OUT STD_LOGIC_VECTOR(0 TO 4);
    Trace_MSR_Reg : OUT STD_LOGIC_VECTOR(0 TO 14);
    Trace_New_Reg_Value : OUT STD_LOGIC_VECTOR(0 TO 31);
    Trace_Jump_Taken : OUT STD_LOGIC;
    Trace_Delay_Slot : OUT STD_LOGIC;
    Trace_Data_Address : OUT STD_LOGIC_VECTOR(0 TO 31);
    Trace_Data_Access : OUT STD_LOGIC;
    Trace_Data_Read : OUT STD_LOGIC;
    Trace_Data_Write : OUT STD_LOGIC;
    Trace_Data_Write_Value : OUT STD_LOGIC_VECTOR(0 TO 31);
    Trace_Data_Byte_Enable : OUT STD_LOGIC_VECTOR(0 TO 3);
    Trace_MB_Halted : OUT STD_LOGIC
  );
END COMPONENT;

-- chipscope 
component trace_icon
  PORT (
    CONTROL0 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CONTROL1 : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0)
	 );
end component;

component trace_ila
  PORT (
    CONTROL : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CLK : IN STD_LOGIC;
    TRIG0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    TRIG1 : IN STD_LOGIC_VECTOR(33 DOWNTO 0);
    TRIG2 : IN STD_LOGIC_VECTOR(8 DOWNTO 0)
	 );
end component;

component trace_vio
  PORT (
    CONTROL : INOUT STD_LOGIC_VECTOR(35 DOWNTO 0);
    CLK : IN STD_LOGIC;
    ASYNC_OUT : OUT STD_LOGIC_VECTOR(1 downto 0);
    SYNC_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));

end component;

-- signals ------------
signal CS_CONTROL0 :  STD_LOGIC_VECTOR(35 DOWNTO 0);
signal CS_CONTROL1 :  STD_LOGIC_VECTOR(35 DOWNTO 0);
signal CS_TRIG0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal CS_TRIG1 :  STD_LOGIC_VECTOR(33 DOWNTO 0);
signal CS_TRIG2 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
signal CS_VIO0 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
signal CS_VIO1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
signal cs_rst: std_logic;
signal cs_stop: std_logic;

-- address range
constant addrBits: integer := 4;
subtype ADDR is std_logic_vector(addrBits - 1 downto 0);

constant idReg: integer := 0;
constant ctlReg: integer := 1;
constant statReg: integer := 2;
constant miscReg: integer := 3;
constant cxReg: integer := 4; -- mandelbrot cx
constant cyReg: integer := 5; -- mandelbrot cy
constant cnReg: integer := 6; -- mandelbrot cy
constant crReg: integer := 7; -- mandelbrot result
constant cxgenMinReg:    integer := 8;  -- cxgen cx_min
constant cxgenDxReg:     integer := 9;  -- cxgen dx
constant cxgenEnableReg: integer := 10; -- cxgen enable
constant cxgenClearReg:  integer := 11; -- cxgen clear
constant mbpipeClearReg: integer := 12; -- mbrot_pipe clear
constant mbpipeCyReg:    integer := 13; -- mbrot_pipe cy
constant startAddrReg:   integer := 14; -- start addr for fr_buff
constant validOutReg:    integer := 15;

constant idAddr:   ADDR :=  std_logic_vector(to_unsigned(idReg,addrBits));
constant ctlAddr:  ADDR :=  std_logic_vector(to_unsigned(ctlReg,addrBits));
constant statAddr: ADDR :=  std_logic_vector(to_unsigned(statReg,addrBits));
constant miscAddr: ADDR :=  std_logic_vector(to_unsigned(miscReg,addrBits));
constant cxAddr: ADDR   :=  std_logic_vector(to_unsigned(cxReg,addrBits));
constant cyAddr: ADDR   :=  std_logic_vector(to_unsigned(cyReg,addrBits));
constant cnAddr: ADDR   :=  std_logic_vector(to_unsigned(cnReg,addrBits));
constant crAddr: ADDR   :=  std_logic_vector(to_unsigned(crReg,addrBits));
constant cxgenMinAddr:    ADDR := std_logic_vector(to_unsigned(cxgenMinReg,addrBits));
constant cxgenDxAddr:     ADDR := std_logic_vector(to_unsigned(cxgenDxReg,addrBits));
constant cxgenEnableAddr: ADDR := std_logic_vector(to_unsigned(cxgenEnableReg,addrBits));
constant cxgenClearAddr:  ADDR := std_logic_vector(to_unsigned(cxgenClearReg,addrBits));
constant mbpipeClearAddr: ADDR := std_logic_vector(to_unsigned(mbpipeClearReg,addrBits));
constant mbpipeCyAddr:    ADDR := std_logic_vector(to_unsigned(mbpipeCyReg,addrBits));
constant startAddr: 		  ADDR := std_logic_vector(to_unsigned(startAddrReg,addrBits)); 
constant validOutAddr:    ADDR := std_logic_vector(to_unsigned(startAddrReg,addrBits)); 

constant ramSelectAddrBit: integer := 29;

-- register set 
type regSet is array(2**addrBits - 1 downto 0) of std_logic_vector(31 downto 0);
signal regs: regSet := (
	idReg => X"00000004",  -- design id
	statReg => X"01020304", 
	cnReg => X"00000020", 
	others => X"00000000");

signal reg_Read_Data: std_logic_vector(31 downto 0);


-- basic core signals
signal IO_Addr_Strobe :  STD_LOGIC;
signal IO_Read_Strobe :  STD_LOGIC;
signal IO_Write_Strobe :  STD_LOGIC;
signal IO_Byte_Address :  STD_LOGIC_VECTOR(31 DOWNTO 0);  -- full address 
signal IO_Address :  STD_LOGIC_VECTOR(addrBits - 1 DOWNTO 0);  -- effective word address 
signal IO_Byte_Enable :  STD_LOGIC_VECTOR(3 DOWNTO 0);
signal IO_Write_Data :  STD_LOGIC_VECTOR(31 DOWNTO 0);
signal IO_Read_Data :  STD_LOGIC_VECTOR(31 DOWNTO 0);
signal IO_Ready :  STD_LOGIC;
signal UART_Interrupt :  STD_LOGIC;
signal FIT1_Interrupt :  STD_LOGIC;
signal FIT2_Interrupt :  STD_LOGIC;
signal PIT1_Interrupt :  STD_LOGIC;
signal PIT2_Interrupt :  STD_LOGIC;
signal GPI1_Interrupt :  STD_LOGIC;
signal GPI2_Interrupt :  STD_LOGIC;
signal INTC_Interrupt :  STD_LOGIC_VECTOR(3 DOWNTO 0);

signal FIT1_Toggle :  STD_LOGIC;
signal PIT1_Toggle :  STD_LOGIC;
signal FIT2_Toggle :  STD_LOGIC;
signal PIT2_Toggle :  STD_LOGIC;
signal PIT2_Enable :  STD_LOGIC;
signal EXT_Interrupt :  STD_LOGIC_VECTOR(2 DOWNTO 0) := (others => '0');
signal INTC_IRQ :  STD_LOGIC;

signal GPO1_i :  STD_LOGIC_VECTOR(7 DOWNTO 0);
signal GPO1_r :  STD_LOGIC_VECTOR(7 DOWNTO 0);  -- pipeline register
signal GPI1_r :  STD_LOGIC_VECTOR(7 DOWNTO 0);  -- pipeline register
signal GPI2_r :  STD_LOGIC_VECTOR(4 DOWNTO 0);  -- pipeline register


-- reset
signal reset: std_logic := '1';  -- general reset
signal areset: std_logic := '1';  -- needed for memory calibration

-- additional logic

signal wrRdy, rdRdy: std_logic;
signal memRdRdy: std_logic := '1' ;

-- simulation bit
signal simStat: std_logic;

-- tracing
signal Trace_PC : STD_LOGIC_VECTOR(0 TO 31);
signal Trace_Instruction : STD_LOGIC_VECTOR(0 TO 31);
signal Trace_Valid_Instr : STD_LOGIC;
signal Trace_Jump_Taken : STD_LOGIC;

signal memPll_ce_0, memPll_ce_90, memPll_lock: std_logic;
signal clkDrp, clk125, clkMem2x, clkMem2x180: std_logic;
signal sysClk, cpuClk: std_logic;
signal stopClk: std_logic := '0';


------------------ memory interface -------------------------
--component dp_mem_wrapper
component dp_mem_wrapper300
--component dp_mem_wrapper250
	generic
	  (
		C3_P0_MASK_SIZE           : integer := 4;
		C3_P0_DATA_PORT_SIZE      : integer := 32;
		C3_P1_MASK_SIZE           : integer := 4;
		C3_P1_DATA_PORT_SIZE      : integer := 32;
		C3_MEMCLK_PERIOD        : integer := 4000; 
											-- Memory data transfer clock period.
		C3_RST_ACT_LOW          : integer := 0; 
											-- # = 1 for active low reset,
											-- # = 0 for active high reset.
		C3_INPUT_CLK_TYPE       : string := "SINGLE_ENDED"; 
											-- input clock type DIFFERENTIAL or SINGLE_ENDED.
		C3_CALIB_SOFT_IP        : string := "TRUE"; 
											-- # = TRUE, Enables the soft calibration logic,
											-- # = FALSE, Disables the soft calibration logic.
		C3_SIMULATION           : string := "FALSE"; 
											-- # = TRUE, Simulating the design. Useful to reduce the simulation time,
											-- # = FALSE, Implementing the design.
		DEBUG_EN                : integer := 0; 
											-- # = 1, Enable debug signals/controls,
											--   = 0, Disable debug signals/controls.
		C3_MEM_ADDR_ORDER       : string := "ROW_BANK_COLUMN"; 
											-- The order in which user address is provided to the memory controller,
											-- ROW_BANK_COLUMN or BANK_ROW_COLUMN.
		C3_NUM_DQ_PINS          : integer := 16; 
											-- External memory data width.
		C3_MEM_ADDR_WIDTH       : integer := 13; 
											-- External memory address width.
		C3_MEM_BANKADDR_WIDTH   : integer := 3 
											-- External memory bank address width.
	  );
  port
  (
	
   mcb_drp_clk                            : in  std_logic;
	async_rst                              : in  std_logic;
	sysclk_2x                              : in  std_logic;
	sysclk_2x_180                          : in  std_logic;
	pll_ce_0                               : in  std_logic;
	pll_ce_90                              : in  std_logic;
	pll_lock                               : in  std_logic;
   calib_done          							: out std_logic;

   mcb3_dram_dq                            : inout  std_logic_vector(15 downto 0);
   mcb3_dram_a                             : out std_logic_vector(12 downto 0);
   mcb3_dram_ba                            : out std_logic_vector(2 downto 0);
   mcb3_dram_ras_n                         : out std_logic;
   mcb3_dram_cas_n                         : out std_logic;
   mcb3_dram_we_n                          : out std_logic;
   mcb3_dram_odt                           : out std_logic;
   mcb3_dram_cke                           : out std_logic;
   mcb3_dram_dm                            : out std_logic;
   mcb3_dram_udqs                          : inout  std_logic;
   mcb3_dram_udqs_n                        : inout  std_logic;
   mcb3_rzq                                : inout  std_logic;
   mcb3_zio                                : inout  std_logic;
   mcb3_dram_udm                           : out std_logic;
   mcb3_dram_dqs                           : inout  std_logic;
   mcb3_dram_dqs_n                         : inout  std_logic;
   mcb3_dram_ck                            : out std_logic;
   mcb3_dram_ck_n                          : out std_logic;
	
	p2_cmd_clk                            : in std_logic;
	p2_cmd_en                             : in std_logic;
	p2_cmd_instr                          : in std_logic_vector(2 downto 0);
	p2_cmd_bl                             : in std_logic_vector(5 downto 0);
	p2_cmd_byte_addr                      : in std_logic_vector(29 downto 0);
	p2_cmd_empty                          : out std_logic;
	p2_cmd_full                           : out std_logic;
	p2_wr_clk                             : in std_logic;
	p2_wr_en                              : in std_logic;
	p2_wr_mask                            : in std_logic_vector(3 downto 0);
	p2_wr_data                            : in std_logic_vector(31 downto 0);
	p2_wr_full                            : out std_logic;
	p2_wr_empty                           : out std_logic;
	p2_wr_count                           : out std_logic_vector(6 downto 0);
	p2_wr_underrun                        : out std_logic;
	p2_wr_error                           : out std_logic;
	p3_cmd_clk                            : in std_logic;
	p3_cmd_en                             : in std_logic;
	p3_cmd_instr                          : in std_logic_vector(2 downto 0);
	p3_cmd_bl                             : in std_logic_vector(5 downto 0);
	p3_cmd_byte_addr                      : in std_logic_vector(29 downto 0);
	p3_cmd_empty                          : out std_logic;
	p3_cmd_full                           : out std_logic;
	p3_rd_clk                             : in std_logic;
	p3_rd_en                              : in std_logic;
	p3_rd_data                            : out std_logic_vector(31 downto 0);
	p3_rd_full                            : out std_logic;
	p3_rd_empty                           : out std_logic;
	p3_rd_count                           : out std_logic_vector(6 downto 0);
	p3_rd_overflow                        : out std_logic;
	p3_rd_error                           : out std_logic;
	p4_cmd_clk                            : in std_logic;
	p4_cmd_en                             : in std_logic;
	p4_cmd_instr                          : in std_logic_vector(2 downto 0);
	p4_cmd_bl                             : in std_logic_vector(5 downto 0);
	p4_cmd_byte_addr                      : in std_logic_vector(29 downto 0);
	p4_cmd_empty                          : out std_logic;
	p4_cmd_full                           : out std_logic;
	p4_wr_clk                             : in std_logic;
	p4_wr_en                              : in std_logic;
	p4_wr_mask                            : in std_logic_vector(3 downto 0);
	p4_wr_data                            : in std_logic_vector(31 downto 0);
	p4_wr_full                            : out std_logic;
	p4_wr_empty                           : out std_logic;
	p4_wr_count                           : out std_logic_vector(6 downto 0);
	p4_wr_underrun                        : out std_logic;
	p4_wr_error                           : out std_logic;
	p5_cmd_clk                            : in std_logic;
	p5_cmd_en                             : in std_logic;
	p5_cmd_instr                          : in std_logic_vector(2 downto 0);
	p5_cmd_bl                             : in std_logic_vector(5 downto 0);
	p5_cmd_byte_addr                      : in std_logic_vector(29 downto 0);
	p5_cmd_empty                          : out std_logic;
	p5_cmd_full                           : out std_logic;
	p5_rd_clk                             : in std_logic;
	p5_rd_en                              : in std_logic;
	p5_rd_data                            : out std_logic_vector(31 downto 0);
	p5_rd_full                            : out std_logic;
	p5_rd_empty                           : out std_logic;
	p5_rd_count                           : out std_logic_vector(6 downto 0);
	p5_rd_overflow                        : out std_logic;
	p5_rd_error                           : out std_logic
  );
end component;

  function getSimString(sim:integer) return string is
  begin
	if sim = 0 then 
		return ("FALSE");
	else 
		return ("TRUE");
	end if;
  end function;
	
  
  signal  calib_done                            : std_logic;

  signal  c3_p2_cmd_en                             : std_logic := '0';
  signal  c3_p2_cmd_instr                          : std_logic_vector(2 downto 0) := (others => '0');
  signal  c3_p2_cmd_bl                             : std_logic_vector(5 downto 0) := (others => '0');
  signal  c3_p2_cmd_byte_addr                      : std_logic_vector(29 downto 0) := (others => '0');
  signal  c3_p2_cmd_empty                          : std_logic;
  signal  c3_p2_cmd_full                           : std_logic;
  signal  c3_p2_wr_en                              : std_logic := '0';
  signal  c3_p2_wr_mask                            : std_logic_vector(3 downto 0) := (others => '0');
  signal  c3_p2_wr_data                            : std_logic_vector(31 downto 0) := (others => '0');
  signal  c3_p2_wr_full                            : std_logic;
  signal  c3_p2_wr_empty                           : std_logic;
  signal  c3_p2_wr_count                           : std_logic_vector(6 downto 0);
  signal  c3_p2_wr_underrun                        : std_logic;
  signal  c3_p2_wr_error                           : std_logic;

  signal  c3_p3_cmd_en                             : std_logic := '0';
  signal  c3_p3_cmd_instr                          : std_logic_vector(2 downto 0) := (others => '0');
  signal  c3_p3_cmd_bl                             : std_logic_vector(5 downto 0) := (others => '0');
  signal  c3_p3_cmd_byte_addr                      : std_logic_vector(29 downto 0) := (others => '0');
  signal  c3_p3_cmd_empty                          : std_logic;
  signal  c3_p3_cmd_full                           : std_logic;
  signal  c3_p3_rd_en                              : std_logic := '0';
  signal  c3_p3_rd_data                            : std_logic_vector(31 downto 0);
  signal  c3_p3_rd_full                            : std_logic;
  signal  c3_p3_rd_empty                           : std_logic;
  signal  c3_p3_rd_count                           : std_logic_vector(6 downto 0);
  signal  c3_p3_rd_overflow                        : std_logic;
  signal  c3_p3_rd_error                           : std_logic;

  signal  c3_p4_cmd_en                             : std_logic := '0';
  signal  c3_p4_cmd_instr                          : std_logic_vector(2 downto 0) := (others => '0');
  signal  c3_p4_cmd_bl                             : std_logic_vector(5 downto 0) := (others => '0');
  signal  c3_p4_cmd_byte_addr                      : std_logic_vector(29 downto 0) := (others => '0');
  signal  c3_p4_cmd_empty                          : std_logic;
  signal  c3_p4_cmd_full                           : std_logic;
  signal  c3_p4_wr_en                              : std_logic := '0';
  signal  c3_p4_wr_mask                            : std_logic_vector(3 downto 0) := (others => '0');
  signal  c3_p4_wr_data                            : std_logic_vector(31 downto 0) := (others => '0');
  signal  c3_p4_wr_full                            : std_logic;
  signal  c3_p4_wr_empty                           : std_logic;
  signal  c3_p4_wr_count                           : std_logic_vector(6 downto 0);
  signal  c3_p4_wr_underrun                        : std_logic;
  signal  c3_p4_wr_error                           : std_logic;

  signal  c3_p5_cmd_en                             : std_logic := '0';
  signal  c3_p5_cmd_instr                          : std_logic_vector(2 downto 0) := (others => '0');
  signal  c3_p5_cmd_bl                             : std_logic_vector(5 downto 0) := (others => '0');
  signal  c3_p5_cmd_byte_addr                      : std_logic_vector(29 downto 0) := (others => '0');
  signal  c3_p5_cmd_empty                          : std_logic;
  signal  c3_p5_cmd_full                           : std_logic;
  signal  c3_p5_rd_en                              : std_logic := '0';
  signal  c3_p5_rd_data                            : std_logic_vector(31 downto 0);
  signal  c3_p5_rd_full                            : std_logic;
  signal  c3_p5_rd_empty                           : std_logic;
  signal  c3_p5_rd_count                           : std_logic_vector(6 downto 0);
  signal  c3_p5_rd_overflow                        : std_logic;
  signal  c3_p5_rd_error                           : std_logic;

  constant single_wr_instr_code: std_logic_vector(2 downto 0) := "000";
  constant burst_wr_instr_code: std_logic_vector(2 downto 0) := "001";
  constant single_rd_instr_code: std_logic_vector(2 downto 0) := "011";
  constant burst_rd_instr_code: std_logic_vector(2 downto 0) := "010";
  constant cpu_bl: std_logic_vector(5 downto 0) := "000000";  -- actual number is 1 more
  constant cpu_wr_mask: std_logic_vector(3 downto 0) := "0000";

  signal cpu_wr_ram_data: std_logic;
  signal cpu_wr_ram_instr: std_logic;
  signal cpu_rd_ram_data: std_logic;
  signal cpu_rd_ram_instr: std_logic;
  signal cpu_ram_addr: std_logic_vector(29 downto 0); -- byte address
  
  signal cxgen_cx_min: std_logic_vector(31 downto 0);
  signal cxgen_dx: std_logic_vector(31 downto 0);
  signal cxgen_enable: std_logic;
  signal cxgen_clear: std_logic;
  signal cxgen_valid: std_logic;
  signal cxgen_cx: std_logic_vector(31 downto 0);
  
  signal mbpipe_clear:     STD_LOGIC;
  signal mbpipe_cy:        STD_LOGIC_VECTOR (31 downto 0);
  signal mbpipe_zx:        STD_LOGIC_VECTOR (31 downto 0);
  signal mbpipe_zy:        STD_LOGIC_VECTOR (31 downto 0);
  signal mbpipe_valid_out: STD_LOGIC;
  signal mbpipe_compare:   STD_LOGIC_VECTOR ((num_mbpipe_stages-1) downto 0);
  
  signal spOColor:         STD_LOGIC_VECTOR(3 downto 0);
  signal spOValid:         STD_LOGIC;
  
  signal colorConverterColorOut: STD_LOGIC_VECTOR (23 downto 0);
  signal colorConverterValidOut: std_logic;

-------------------------------------------------------------
component cxgen is
    Port ( cx_min : in  STD_LOGIC_VECTOR (31 downto 0);
           dx     : in  STD_LOGIC_VECTOR (31 downto 0);
           enable : in  STD_LOGIC;
           clear  : in  STD_LOGIC;
           reset  : in  STD_LOGIC;
           clk    : in  STD_LOGIC;
           cx     : out STD_LOGIC_VECTOR (31 downto 0);
           valid  : out STD_LOGIC);
end component;

-------------------------------------------------------------

component mbrot_pipe is
  generic( num_cx     : integer := 800;
           num_stages : integer := 16);
    Port ( clk        : in   STD_LOGIC;
           reset      : in   STD_LOGIC;
           clear      : in   STD_LOGIC;
           valid_in   : in   STD_LOGIC;
           cx         : in   STD_LOGIC_VECTOR (31 downto 0);
           cy         : in   STD_LOGIC_VECTOR (31 downto 0);
           zx         : out  STD_LOGIC_VECTOR (31 downto 0);
           zy         : out  STD_LOGIC_VECTOR (31 downto 0);
           valid_out  : out  STD_LOGIC;
           compare    : out  STD_LOGIC_VECTOR ((num_stages-1) downto 0));
end component;

-------------------------------------------------------------
 
COMPONENT shiftPipe
generic (width: integer := 4; depth: integer := 16);
port
(
  clk, reset:	in std_logic;
  iCmpVector:	in std_logic_vector(depth-1 downto 0);
  iValid:		in std_logic;

  oColor:		out std_logic_vector(width-1 downto 0);
  oValid:		out std_logic
);
END COMPONENT;
-------------------------------------------------------------

COMPONENT ColorConverter_4_24 is
    Port ( clock : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           color_in : in  STD_LOGIC_VECTOR (3 downto 0);
           color_out : out  STD_LOGIC_VECTOR (23 downto 0);
           valid_in: in std_logic;
           valid_out: out std_logic);
end COMPONENT;
  
-------------------------------------------------------------
	COMPONENT dp_mem_infrastructure
	  generic (
			hasDram: integer := 1;
			simulation: integer := 0;
			trace: integer := 1  -- use chipscope
	  );
	PORT(
		clkIn : IN std_logic;
		stopCpu : IN std_logic;
		extRstIn_n : IN std_logic;
		intRstIn : IN std_logic;          
		clkSys : OUT std_logic;
		clkCpu : OUT std_logic;
		clk125 : OUT std_logic;
		clkDrp : OUT std_logic;
		clkMem2x : OUT std_logic;
		clkMem2x180 : OUT std_logic;
		memPll_ce_0 : OUT std_logic;
		memPll_ce_90 : OUT std_logic;
		memPll_lock : OUT std_logic;
		areset        : out std_logic;	-- early reset, clocked with input clock
		dreset        : out std_logic	-- delayed, synchronous reset
		);
	END COMPONENT;
-------------------------------------------------------------

	COMPONENT hdmiOutIF
	generic (
		xga: integer := 1; -- xga or 720p on hdmi
		simulation: integer := 0
	);
	PORT(
		CLK100_IN : IN std_logic;
		hdmiDataR : IN std_logic_vector(7 downto 0);
		hdmiDataG : IN std_logic_vector(7 downto 0);
		hdmiDataB : IN std_logic_vector(7 downto 0);
		RESET : IN std_logic;          
		clkHdmiTx : OUT std_logic;
		hdmiHsync	: out std_logic;  -- row sync for address generator
		hdmiVsync	: out std_logic;  -- frame sync for address generator
		hdmiHsyncIn			: in std_logic;  -- row sync from data source
		hdmiVsyncIn			: in std_logic;  -- vsync from data source
		hdmiFsync   : out std_logic;  -- frame sync. active with very last row 
		hdmiActive	: out std_logic;  -- read enable
		hdmiActiveIn	: in std_logic;  -- read enable
		hdmiTx0_p : OUT std_logic;
		hdmiTx0_n : OUT std_logic;
		hdmiTx1_p : OUT std_logic;
		hdmiTx1_n : OUT std_logic;
		hdmiTx2_p : OUT std_logic;
		hdmiTx2_n : OUT std_logic;
		hdmiTx3_p : OUT std_logic;
		hdmiTx3_n : OUT std_logic
	);
	END COMPONENT;

signal clkHdmiTx : std_logic;
signal hdmiDataRTx : std_logic_vector(7 downto 0) := X"55";
signal hdmiDataGTx : std_logic_vector(7 downto 0) := X"11";
signal hdmiDataBTx : std_logic_vector(7 downto 0) := X"F0";
signal hdmiHsyncTx : std_logic;
signal hdmiVsyncTx : std_logic;
signal hdmiHsyncTxIn : std_logic;
signal hdmiVsyncTxIn : std_logic;
signal hdmiFsyncTx : std_logic;
signal hdmiActiveTx :std_logic;
signal hdmiActiveTxIn :std_logic;

signal line_length: integer := 1024;

function getXgaMode return std_logic is
begin
	if xga /= 0 then
		return '1';
	else
		return '0';
	end if;
end function;

-------------------------------------------------------------
COMPONENT dram_reader
  generic (
		xga: integer := 1; -- xga or 720p on hdmi
		simulation: integer := 0
  );
    Port ( 
		clk : in  STD_LOGIC;
		rst : in  STD_LOGIC;
		hsync : in  STD_LOGIC;
		vsync : in  STD_LOGIC;
		fsync : in  STD_LOGIC;
		active : in  STD_LOGIC;
		active_out : out  STD_LOGIC;
		hsync_out : out  STD_LOGIC;
		vsync_out : out  STD_LOGIC;
		cmd : out  STD_LOGIC_VECTOR (2 downto 0);
		cmdEn : out  STD_LOGIC;
		cmdFull : in  STD_LOGIC;
		cmdBl : out  STD_LOGIC_vector(5 downto 0);
		frameBase: std_logic_vector(29 downto 0);
		addr : out  STD_LOGIC_VECTOR (29 downto 0);
		rdEn : out  STD_LOGIC;
		rdEmpty : in  STD_LOGIC;
		rdFull : in  STD_LOGIC;
		rdData : in  STD_LOGIC_VECTOR (31 downto 0);
		data : out  STD_LOGIC_VECTOR (31 downto 0)
	);
END COMPONENT;

signal imageDataTx: std_logic_vector(31 downto 0);
constant frameBase: std_logic_vector(29 downto 0) := (others => '0');
constant frame2Base: std_logic_vector(29 downto 0) := (22 => '1', others => '0');
signal frameBaseTx: std_logic_vector(29 downto 0);
signal frameBaseRx: std_logic_vector(29 downto 0);
signal hdmiReset: std_logic;
signal vsyncTx: std_logic;
signal hsyncTx: std_logic;
signal activeTx: std_logic;

-------------------------------------------------------------
    COMPONENT mbrot
	 generic (maxDsp: integer := 1; latency: integer := 3);
    PORT(
         cx : IN  std_logic_vector(31 downto 0);
         cy : IN  std_logic_vector(31 downto 0);
         nmax : IN  std_logic_vector(31 downto 0);
         n : OUT  std_logic_vector(31 downto 0);
         done : OUT  std_logic;
         clk : IN  std_logic;
         rst : IN  std_logic
        );
    END COMPONENT;

signal mb_n, mb_n_i: std_logic_vector(31 downto 0);
signal mb_rst: std_logic; -- write pulse on cx register
signal mb_done, mb_done_i: std_logic; 

signal cxReg_i :  std_logic_vector(31 downto 0);
signal cyReg_i :  std_logic_vector(31 downto 0);
signal cnReg_i :  std_logic_vector(31 downto 0);

-------------------------------------------------------------
	COMPONENT hdmiRx
	PORT(
		hdmiRx_p : IN std_logic_vector(3 downto 0);
		hdmiRx_n : IN std_logic_vector(3 downto 0);
		reset : IN std_logic;          
		pclk : OUT std_logic;
		frame_width     : OUT std_logic_vector(15 downto 0) := (others => '0');
		frame_height    : OUT std_logic_vector(15 downto 0) := (others => '0');
		new_frame     : OUT std_logic;
		line_end     : OUT std_logic;
		hsync : OUT std_logic;
		vsync : OUT std_logic;
		de : OUT std_logic;
		red : OUT std_logic_vector(7 downto 0);
		green : OUT std_logic_vector(7 downto 0);
		blue : OUT std_logic_vector(7 downto 0)
		);
	END COMPONENT;

signal clkHdmiRx : std_logic;
	
signal hdmiRxClk: std_logic;
signal hdmiRxHsync: std_logic;
signal hdmiRxVsync: std_logic;
signal hdmiRxActive: std_logic;
signal hdmiRxRed: std_logic_vector(7 downto 0);
signal hdmiRxGreen: std_logic_vector(7 downto 0);
signal hdmiRxBlue: std_logic_vector(7 downto 0);
signal hdmiRx_new_frame     : std_logic;
signal hdmiRx_line_end     : std_logic;
signal hdmiRx_frame_width     : std_logic_vector(15 downto 0) := (others => '0');
signal hdmiRx_frame_height    : std_logic_vector(15 downto 0) := (others => '0');

signal hdmiRxDreg0, hdmiRxDreg1: std_logic_vector(23 downto 0);
signal hdmiRxAct_r0, hdmiRxAct_r1: std_logic;

-------------------------------------------------------------
-- hdmi edid
COMPONENT i2cSlave
PORT(
	clk : IN std_logic;
	rst : IN std_logic;
	scl : IN std_logic;       
	sda : INOUT std_logic
	);
END COMPONENT;

-------------------------------------------------------------

begin

  -- simulation mode detection
  simMode: if simulation /= 0 generate
  begin
	simStat <= '1';
  end generate;
  impMode: if simulation = 0 generate
  begin
	simStat <= '0';
  end generate;
  
  -- cxgen
  cxgen_cx_min <= regs(cxgenMinReg);
  cxgen_dx     <= regs(cxgenDxReg);
  cxgen_enable <= regs(cxgenEnableReg)(0);
  cxgen_clear  <= regs(cxgenClearReg)(0);
  CXGEN_I: cxgen port map (
    cx_min => cxgen_cx_min,
	  dx     => cxgen_dx,
	  enable => cxgen_enable,
	  clear  => cxgen_clear,
	  reset  => reset,
	  clk    => clk,
	  cx     => cxgen_cx,
	  valid  => cxgen_valid
  );
 
  -- mbrot_pipe
  mbpipe_cy    <= regs(mbpipeCyReg);
  mbpipe_clear <= regs(mbpipeClearReg)(0);
  MBPIPE_I: mbrot_pipe
    generic map (num_cx     => num_cx,
                 num_stages => num_mbpipe_stages)
    port map    (clk       => clk,
                 reset     => reset,
                 clear     => mbpipe_clear,
                 valid_in  => cxgen_valid,
                 cx        => cxgen_cx,
                 cy        => mbpipe_cy,
                 zx        => mbpipe_zx,
                 zy        => mbpipe_zy,
                 valid_out => mbpipe_valid_out,
                 compare   => mbpipe_compare
  );
  
  -- shiftPipe
   SHIFTPIPE_I: shiftPipe
   generic map (width => 4, depth => num_mbpipe_stages)
   PORT MAP (
          clk => clk,
          reset => reset,
          iCmpVector => mbpipe_compare,
          iValid => mbpipe_valid_out,
          oColor => spOColor,
          oValid => spOValid
        );
       
  -- ColorConverter
  COLERCONVERTER_I: ColorConverter_4_24 port map (
    clock => clk,
    reset => reset,
    color_in => spOColor,
    color_out => colorConverterColorOut,
    valid_in => spOValid,
    valid_out => colorConverterValidOut);

  -- infrastructure: clock and reset
	clkRst: dp_mem_infrastructure PORT MAP(
		clkIn => clk,
		clkSys => sysClk,
		stopCpu => stopClk,
		clkCpu => cpuClk,
		clk125 => clk125,
		clkDrp => clkDrp,
		clkMem2x => clkMem2x,
		clkMem2x180 => clkMem2x180,
		memPll_ce_0 => memPll_ce_0,
		memPll_ce_90 => memPll_ce_90,
		memPll_lock => memPll_lock,
		extRstIn_n => rst_n,
		intRstIn => cs_rst,
		areset => areset, -- reset for dram only
		dreset => reset
	);
  
	-------------------------------
	-------------------------------
	-- use the instance name as given in xco file. Otherwise edit .bmm file 
	
  mcs_0 : mblaze
  PORT MAP (
	 Clk => cpuClk,
	 Reset => Reset,
	 IO_Addr_Strobe => IO_Addr_Strobe,
	 IO_Read_Strobe => IO_Read_Strobe,
	 IO_Write_Strobe => IO_Write_Strobe,
	 IO_Address => IO_Byte_Address,
	 IO_Byte_Enable => IO_Byte_Enable,
	 IO_Write_Data => IO_Write_Data,
	 IO_Read_Data => IO_Read_Data,
	 IO_Ready => IO_Ready,
	 UART_Rx => UART_Rx,
	 UART_Tx => UART_Tx,
	 UART_Interrupt => UART_Interrupt,
	 FIT1_Interrupt => FIT1_Interrupt,
	 FIT1_Toggle => FIT1_Toggle,
	 FIT2_Interrupt => FIT2_Interrupt,
	 FIT2_Toggle => FIT2_Toggle,
	 PIT1_Interrupt => PIT1_Interrupt,
	 PIT1_Toggle => PIT1_Toggle,
	 PIT2_Enable => PIT2_Enable,
	 PIT2_Interrupt => PIT2_Interrupt,
	 PIT2_Toggle => PIT2_Toggle,
	 GPO1 => GPO1_i,
	 GPI1 => GPI1_r,
	 GPI2 => GPI2_r,
	 GPI1_Interrupt => GPI1_Interrupt,
	 GPI2_Interrupt => GPI2_Interrupt,
	 INTC_Interrupt => EXT_Interrupt,
	 INTC_IRQ => INTC_IRQ,
	 Trace_Instruction => Trace_Instruction,
	 Trace_Valid_Instr => Trace_Valid_Instr,
	 Trace_Jump_Taken => Trace_Jump_Taken,
	 Trace_PC => Trace_PC
  );

	-- with trace enabled, we can add logic to set HW breakpoints and stop the clock
	withTrace: if trace /= 0 generate
	begin
		
		-- insert chipscope if not in simulation mode
		-- no chipscope
		withChipscope: if false generate -- simulation = 0 generate
		begin

			csCtl : trace_icon
			  port map (
				 CONTROL0 => CS_CONTROL0,
				 CONTROL1 => CS_CONTROL1
				 );
			csIla : trace_ila
			  port map (
				 CONTROL => CS_CONTROL0,
				 CLK => sysClk,
				 TRIG0 => CS_TRIG0,
				 TRIG1 => CS_TRIG1,
				 TRIG2 => CS_TRIG2
				 );
			
			-- registered map
			process
			begin
			wait until rising_edge(sysClk);
				cs_trig0 <= Trace_PC;
				cs_trig1 <= Trace_Instruction & Trace_Valid_Instr & Trace_Jump_Taken;
				CS_TRIG2(7 downto 0) <= EXT_Interrupt & UART_Interrupt & FIT1_Interrupt & FIT2_Interrupt & PIT1_Interrupt & PIT2_Interrupt;
				cs_trig2(8) <= INTC_IRQ;
			end process;
			
			csVio : trace_vio
			  port map (
				 CONTROL => CS_CONTROL1,
				 CLK => sysClk,
				 ASYNC_OUT => CS_VIO0,
				 SYNC_OUT => CS_VIO1);
				 
			-- registered map
			process
			begin
			wait until rising_edge(sysClk);
				cs_rst <= CS_VIO0(0);
				-- stop on address match
				if (cs_vio0(1) = '1') and (CS_VIO1 = Trace_PC) then
					cs_stop <= '1';
				else
					cs_stop <= '0';
				end if;
			end process;

		end generate;
		
		noChipscope: if simulation /= 0 generate
		begin
			cs_rst <= '0';	-- force reset to 0
			cs_stop <= '0';
		end generate;

		-- no other action at the moment
		stopClk <= cs_stop; 
	end generate;
	
  -- effective address
  IO_Address <= IO_Byte_Address(addrBits + 1 downto 2); -- make word address
  
  -- ready logic
  IO_Ready <= wrRdy or rdRdy;
  

  -- write control
  wrProc: process
  begin
		wait until rising_edge(cpuClk);
		if reset = '1' then
			regs(ctlReg) <= (others => '0');
			regs(miscReg) <= (others => '0');
		else
			if IO_Write_Strobe = '1' then
				wrRdy <= '1';
				
				if (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = ctlAddr) then
					regs(ctlreg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = miscAddr) then
					regs(miscReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cxAddr) then
					regs(cxReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cyAddr) then
					regs(cyReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cnAddr) then
					regs(cnReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cxgenMinAddr) then
					regs(cxgenMinReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cxgenDxAddr) then
					regs(cxgenDxReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cxgenEnableAddr) then
					regs(cxgenEnableReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = cxgenClearAddr) then
					regs(cxgenClearReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = mbpipeClearAddr) then
					regs(mbpipeClearReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = mbpipeCyAddr) then
					regs(mbpipeCyReg) <= IO_Write_Data;
				elsif (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0) = startAddr) then
					regs(startAddrReg) <= IO_Write_Data;
				end if;
				
			else
				wrRdy <= '0';
			end if;
		end if;
  end process;
  
  -- status map
  statMap: block
  begin
		 regs(statReg)(31) <= simStat;
		 regs(statReg)(30) <= FIT1_Toggle;
		 regs(statReg)(29) <= INTC_IRQ;
		 regs(statReg)(28) <= calib_done;
		 
		 regs(statReg)(27) <= c3_p2_cmd_empty;
		 regs(statReg)(26) <= c3_p2_cmd_full;
		 regs(statReg)(25) <= c3_p2_wr_empty;
		 regs(statReg)(24) <= c3_p2_wr_full;
		 regs(statReg)(23) <= c3_p3_cmd_empty;
		 regs(statReg)(22) <= c3_p3_cmd_full;
		 regs(statReg)(21) <= c3_p3_rd_empty;
		 regs(statReg)(20) <= c3_p3_rd_full;

		 regs(statReg)(19) <= getXgaMode;
		 
		 regs(statReg)(18) <= mb_done;

		 regs(statReg)(17 downto 0) <= (others => '0');
  end block;

  -- control map
  ctlMap: block
  begin
		EXT_Interrupt <= regs(ctlReg)(5 downto 3);
		PIT2_Enable <= regs(ctlReg)(2);
  end block;
  
  -- read control
  rdBlock: block
  begin
		-- data mux
		-- regs
		-- use register address with regs
		with IO_Address(addrBits - 1 downto 0) select
			reg_Read_Data <= regs(idReg) when idAddr,
								 regs(ctlReg) when ctlAddr,
								 regs(statReg) when statAddr,
								 regs(miscReg) when miscAddr,
                 regs(validOutReg) when validOutAddr,
								 mb_n when crAddr,
								 (others => '0') when others;
		-- memory						 
		-- use byte address to select reg vs mem
		with IO_Byte_Address(ramSelectAddrBit) select
			IO_Read_Data <= c3_p3_rd_data when '1', reg_Read_Data when others;
			
		-- ready
		with IO_Byte_Address(ramSelectAddrBit) select
			rdRdy <= memRdRdy when '1', IO_Read_Strobe when others;
			
  end block;
  
  -- input pipeline
  gpinPIpe: process
  begin
		wait until rising_edge(sysClk);
		gpi1_r <= gpi1;
		gpi2_r <= gpi2;
  end process;
  
  -- output pipeline
  gpoutPIpe: process
  begin
		wait until rising_edge(sysClk);
		gpo1 <= gpo1_r;
  end process;

  -- output mux LED vs PI toggle 
  ledMux: block
  begin
		gpo1_r(7 downto 2) <= gpo1_i(7 downto 2);
		gpo1_r(1) <= gpo1_i(1) when regs(ctlReg)(1) = '0' else PIT2_Toggle;
		gpo1_r(0) <= gpo1_i(0) when regs(ctlReg)(0) = '0' else PIT1_Toggle;
  end block;
 
  withDram: if hasDram /= 0 generate
  begin

	-- atlys has pulldown on chip_select
	-- mcb3_dram_cs_n <= '0';
	cpu_ram_addr(29 downto ramSelectAddrBit) <= (others => '0');
	cpu_ram_addr(ramSelectAddrBit - 1 downto 2) <= (IO_Byte_Address(ramSelectAddrBit - 1 downto 2));
	cpu_ram_addr(1 downto 0) <= (others => '0');
	
	cpu_rd_ram_instr <= '1' when IO_Read_Strobe = '1' and IO_Byte_Address(ramSelectAddrBit) = '1' else '0';
	-- cpu_rd_ram_data <= '1' when IO_Read_Strobe = '1' and IO_Byte_Address(ramSelectAddrBit) = '1' else '0';
	cpu_wr_ram_data <= '1' when IO_Write_Strobe = '1' and IO_Byte_Address(ramSelectAddrBit) = '1' else '0';

	-- read access waiting for data
	process
		variable wt: std_logic;
	begin
		wait until rising_edge(cpuClk);
		if reset = '1' then 
			wt := '0';
		elsif cpu_rd_ram_instr = '1' then
			wt := '1';
		elsif cpu_rd_ram_data = '1' then
			wt := '0';
		end if;
		
		-- read data access when data available (not empty)
		if wt = '1' and c3_p3_rd_empty = '0' then 
			cpu_rd_ram_data <= '1';
		else
			cpu_rd_ram_data <= '0';
		end if;

	end process;

	-- read ready whith read data
	memRdRdy <= cpu_rd_ram_data;

	
	-- write instruction delayed wrt data write
	process
	begin
		wait until rising_edge(cpuClk);
		cpu_wr_ram_instr <= cpu_wr_ram_data;
	end process;
	
	
--	Inst_dp_mem_wrapper: dp_mem_wrapper
--	Inst_dp_mem_wrapper: dp_mem_wrapper250
	Inst_dp_mem_wrapper: dp_mem_wrapper300 
	generic map ( C3_SIMULATION => getSimString(simulation)) -- C3_SIMULATION)
	PORT MAP (
		mcb3_dram_dq                         => mcb3_dram_dq,
		mcb3_dram_a                          => mcb3_dram_a,
		mcb3_dram_ba                         => mcb3_dram_ba,
		mcb3_dram_ras_n                      => mcb3_dram_ras_n,
		mcb3_dram_cas_n                      => mcb3_dram_cas_n,
		mcb3_dram_we_n                       => mcb3_dram_we_n,
		mcb3_dram_odt                        => mcb3_dram_odt,
		mcb3_dram_cke                        => mcb3_dram_cke,
		mcb3_dram_dm                         => mcb3_dram_dm,
		mcb3_dram_udqs                       => mcb3_dram_udqs,
		mcb3_dram_udqs_n                     => mcb3_dram_udqs_n,
		mcb3_rzq                             => mcb3_rzq,
		mcb3_zio                             => mcb3_zio,
		mcb3_dram_udm                        => mcb3_dram_udm,
		mcb_drp_clk                    		 => clkDrp,
		mcb3_dram_dqs                        => mcb3_dram_dqs,
		mcb3_dram_dqs_n                      => mcb3_dram_dqs_n,
		mcb3_dram_ck                         => mcb3_dram_ck,
		mcb3_dram_ck_n                       => mcb3_dram_ck_n,
		-- 
		p2_cmd_clk                           =>  cpuClk,
		p2_cmd_en                            =>  cpu_wr_ram_instr,
		p2_cmd_instr                         =>  single_wr_instr_code,
		p2_cmd_bl                            =>  cpu_bl,
		p2_cmd_byte_addr                     =>  cpu_ram_addr,
		p2_cmd_empty                         =>  c3_p2_cmd_empty,
		p2_cmd_full                          =>  c3_p2_cmd_full,
		p2_wr_clk                            =>  cpuClk,
		p2_wr_en                             =>  cpu_wr_ram_data,
		p2_wr_mask                           =>  cpu_wr_mask,
		p2_wr_data                           =>  IO_Write_Data,
		p2_wr_full                           =>  c3_p2_wr_full,
		p2_wr_empty                          =>  c3_p2_wr_empty,
		p2_wr_count                          =>  c3_p2_wr_count,
		p2_wr_underrun                       =>  c3_p2_wr_underrun,
		p2_wr_error                          =>  c3_p2_wr_error,
		
		p3_cmd_clk                           =>  cpuClk,
		p3_cmd_en                            =>  cpu_rd_ram_instr,
		p3_cmd_instr                         =>  single_rd_instr_code,
		p3_cmd_bl                            =>  cpu_bl,
		p3_cmd_byte_addr                     =>  cpu_ram_addr,
		p3_cmd_empty                         =>  c3_p3_cmd_empty,
		p3_cmd_full                          =>  c3_p3_cmd_full,
		p3_rd_clk                            =>  cpuClk,
		p3_rd_en                             =>  cpu_rd_ram_data,
		p3_rd_data                           =>  c3_p3_rd_data,
		p3_rd_full                           =>  c3_p3_rd_full,
		p3_rd_empty                          =>  c3_p3_rd_empty,
		p3_rd_count                          =>  c3_p3_rd_count,
		p3_rd_overflow                       =>  c3_p3_rd_overflow,
		p3_rd_error                          =>  c3_p3_rd_error,

		p4_cmd_clk                           =>  clk,
		p4_cmd_en                            =>  c3_p4_cmd_en,
		p4_cmd_instr                         =>  c3_p4_cmd_instr,
		p4_cmd_bl                            =>  c3_p4_cmd_bl,
		p4_cmd_byte_addr                     =>  c3_p4_cmd_byte_addr,
		p4_cmd_empty                         =>  c3_p4_cmd_empty,
		p4_cmd_full                          =>  c3_p4_cmd_full,
		p4_wr_clk                            =>  clk,
		p4_wr_en                             =>  c3_p4_wr_en,
		p4_wr_mask                           =>  c3_p4_wr_mask,
		p4_wr_data                           =>  c3_p4_wr_data,
		p4_wr_full                           =>  c3_p4_wr_full,
		p4_wr_empty                          =>  c3_p4_wr_empty,
		p4_wr_count                          =>  c3_p4_wr_count,
		p4_wr_underrun                       =>  c3_p4_wr_underrun,
		p4_wr_error                          =>  c3_p4_wr_error,

		p5_cmd_clk                           =>  clkHdmiTx,
		p5_cmd_en                            =>  c3_p5_cmd_en,
		p5_cmd_instr                         =>  c3_p5_cmd_instr,
		p5_cmd_bl                            =>  c3_p5_cmd_bl,
		p5_cmd_byte_addr                     =>  c3_p5_cmd_byte_addr,
		p5_cmd_empty                         =>  c3_p5_cmd_empty,
		p5_cmd_full                          =>  c3_p5_cmd_full,
		p5_rd_clk                            =>  clkHdmiTx,
		p5_rd_en                             =>  c3_p5_rd_en,
		p5_rd_data                           =>  c3_p5_rd_data,
		p5_rd_full                           =>  c3_p5_rd_full,
		p5_rd_empty                          =>  c3_p5_rd_empty,
		p5_rd_count                          =>  c3_p5_rd_count,
		p5_rd_overflow                       =>  c3_p5_rd_overflow,
		p5_rd_error                          =>  c3_p5_rd_error,
		--
		calib_done                      => calib_done,
		async_rst                       => areset,  -- memory reset
		sysclk_2x                       => clkMem2x,
		sysclk_2x_180                   => clkMem2x180,
		pll_ce_0                        => memPll_ce_0,
		pll_ce_90                       => memPll_ce_90,
		pll_lock                        => memPll_lock
	);

  
  end generate;  
  
  withHdmiTx: if hasHdmiTx /= 0 generate
  begin
  
		Inst_hdmiOutIF: hdmiOutIF 
		generic map ( xga => xga, simulation => simulation)
		PORT MAP(
			CLK100_IN => sysClk,
			clkHdmiTx => clkHdmiTx,
			hdmiDataR => hdmiDataRTx,
			hdmiDataG => hdmiDataGTx,
			hdmiDataB => hdmiDataBTx,
			hdmiHsync => hdmiHsyncTx,
			hdmiVsync => hdmiVsyncTx,
			hdmiHsyncIn => hdmiHsyncTxIn,
			hdmiVsyncIn => hdmiVsyncTxIn,
			hdmiFsync => hdmiFsyncTx,
			hdmiActive => hdmiActiveTx,
			hdmiActiveIn => hdmiActiveTxIn,
			hdmiTx0_p => hdmiTx0_p,
			hdmiTx0_n => hdmiTx0_n,
			hdmiTx1_p => hdmiTx1_p,
			hdmiTx1_n => hdmiTx1_n,
			hdmiTx2_p => hdmiTx2_p,
			hdmiTx2_n => hdmiTx2_n,
			hdmiTx3_p => hdmiTx3_p,
			hdmiTx3_n => hdmiTx3_n,
			RESET => hdmiReset
		);
	-- test: change color every frame

	frameBaseTx <= frameBase when gpi1(7) = '0' else frame2Base;
	frameBaseRx <= frameBase when gpi1(6) = '1' else frame2Base;

	Inst_dram_reader: dram_reader 
	generic map ( xga => xga, simulation => simulation)
	PORT MAP(
		clk => clkHdmiTx,
		rst => hdmiReset,
		hsync => hdmiHsyncTx,
		vsync => hdmiVsyncTx,
		fsync => hdmiFsyncTx,
		hsync_out => hsyncTx,
		vsync_out => vsyncTx,
		frameBase => frameBaseTx,
		active => hdmiActiveTx,
		active_out => activeTx,
		cmd => c3_p5_cmd_instr,
		cmdEn => c3_p5_cmd_en,
		cmdBl => c3_p5_cmd_bl,
		addr => c3_p5_cmd_byte_addr,
		rdEmpty => c3_p5_rd_empty,
		rdData => c3_p5_rd_data,
		rdEn => c3_p5_rd_en,
		data => imageDataTx,
		cmdFull => c3_p5_cmd_full,
		rdFull => c3_p5_rd_full
	);

	hdmiReset <= reset or not calib_done;
	

	process
		variable greyval: std_logic_vector(7 downto 0);
		constant threshold: std_logic_vector(7 downto 0) := X"5f";
	begin
		wait until rising_edge(clkHdmiTx);
		-- rgb 
		if gpi1(2 downto 0) = "000" then
			hdmiDataBTx <= imageDataTx( 7 downto  0);
			hdmiDataRTx <= imageDataTx(15 downto  8);
			hdmiDataGTx <= imageDataTx(23 downto 16);
			hdmiHsyncTxIn <= hsyncTx;
			hdmiVsyncTxIn <= vsyncTx;
			hdmiActiveTxIn <= activeTx;
		elsif gpi1(2 downto 0) = "001" then
			hdmiDataBTx <= X"F0";
			hdmiDataRTx <= X"55";
			hdmiDataGTx <= X"10";
			hdmiHsyncTxIn <= hdmiHsyncTx;
			hdmiVsyncTxIn <= hdmiVsyncTx;
			hdmiActiveTxIn <= hdmiActiveTx;
		-- grey
		elsif gpi1(2 downto 0) = "010" then
			hdmiDataBTx <= imageDataTx( 7 downto  0);
			hdmiDataRTx <= imageDataTx( 7 downto  0);
			hdmiDataGTx <= imageDataTx( 7 downto  0);
			hdmiHsyncTxIn <= hsyncTx;
			hdmiVsyncTxIn <= vsyncTx;
			hdmiActiveTxIn <= activeTx;
		elsif gpi1(2 downto 0) = "011" then
			hdmiDataBTx <= X"F0";
			hdmiDataRTx <= X"F0";
			hdmiDataGTx <= X"F0";
			hdmiHsyncTxIn <= hdmiHsyncTx;
			hdmiVsyncTxIn <= hdmiVsyncTx;
			hdmiActiveTxIn <= hdmiActiveTx;
		else
			greyval := imageDataTx( 7 downto  0) or imageDataTx(15 downto  8) or imageDataTx(23 downto 16);
			if greyval > threshold then
				hdmiDataBTx <= X"FF";
				hdmiDataRTx <= X"FF";
				hdmiDataGTx <= X"FF";
			else
				hdmiDataBTx <= X"00";
				hdmiDataRTx <= X"00";
				hdmiDataGTx <= X"00";
			end if;
			hdmiHsyncTxIn <= hsyncTx;
			hdmiVsyncTxIn <= vsyncTx;
			hdmiActiveTxIn <= activeTx;
		end if;
	end process;

  end generate;

	withMbrot: if hasMbrot /= 0 generate
	begin
		mb_rst <= '1' when (IO_Write_Strobe = '1') and (IO_Byte_Address(ramSelectAddrBit) = '0') and (IO_Address(addrBits - 1 downto 0)) = cxAddr else '0';
		
		-- input and output pipeline required for speed
		process
		begin
			wait until rising_edge(cpuClk);
			cxReg_i <= regs(cxReg);
			cyReg_i <= regs(cyReg);
			cnReg_i <= regs(cnReg);
			mb_n <= mb_n_i;
			mb_done <= mb_done_i;
		end process;
	
		mbCompute: mbrot 
		generic map (maxDsp => 0, latency => 3) -- maybe we need maxDsp = 1 for 100MHz
		PORT MAP (
		 cx => cxReg_i,
		 cy => cyReg_i,
		 nmax => cnReg_i,
		 n => mb_n_i,
		 done => mb_done_i,
		 clk => cpuClk,
		 rst => mb_rst
	  );

	end generate;
 

		process
			variable cnt : integer range 0 to 32 := 0;
			variable row_base_addr  : std_logic_vector(29 downto 0) := (others => '0');
		begin
			wait until rising_edge(clk);
      
      if hdmiRxActive = '0' then
        cnt := 0;
				c3_p4_cmd_en <= '1';
        c3_p4_cmd_byte_addr <= regs(startAddrReg)(29 downto 0);
      else
				if cnt = 31 then
					cnt := 0;
					c3_p4_cmd_en <= '1';
					c3_p4_cmd_byte_addr <= c3_p4_cmd_byte_addr + 32*4;
				else
					cnt := cnt + 1;
				end if;
      end if;
		end process;

		-- direct write signals
		c3_p4_cmd_instr <= single_wr_instr_code;
		c3_p4_cmd_bl <= std_logic_vector(to_unsigned(31, 6));
		c3_p4_wr_mask <= "0000";
		
		-- pipelined write signals
		process
		begin
			wait until rising_edge(clk);
         regs(validOutReg)(3) <= colorConverterValidOut;
			hdmiRxact_r0 <= colorConverterValidOut;
			hdmiRxact_r1 <= hdmiRxact_r0;
			hdmiRxdreg0  <= colorConverterColorOut;
			hdmiRxdreg1  <= hdmiRxdreg0;
			if (hdmiRxact_r0 = '0') and (hdmiRxact_r1 = '0') then -- supress single cycle actives from rx decoder
				c3_p4_wr_en <= '0';
			elsif (hdmiRxact_r0 = '1') and (hdmiRxact_r1 = '1') then -- supress single cycle actives from rx decoder
				c3_p4_wr_en <= '1';
			elsif (hdmiRxact_r0 = '0') and (hdmiRxact_r1 = '1') and (c3_p4_wr_en = '1')  then
				c3_p4_wr_en <= '1';
			else
				c3_p4_wr_en <= '0';
			end if;

			c3_p4_wr_data <= X"00" & hdmiRxdreg1;
--			if (hdmiRxActive = '1') and (hdmiRxVsync = '0') then -- block 
--				c3_p4_wr_en <= '1';
--			else
--				c3_p4_wr_en <= '0';
--			end if;
--			c3_p4_wr_data <= X"00" & hdmiRxRed & hdmiRxGreen & hdmiRxBlue;
		end process;
 
end rtl;
